module check
pub fn add(x u64, y u64) u64 {
   return x + y
}
